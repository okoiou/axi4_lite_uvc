
package axi4_lite_env_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;
import axi4_lite_pkg::*;
`include "axi4_lite_virtual_sequencer.sv"
`include "axi4_lite_virtual_sequence.sv"
`include "axi4_lite_env_cfg.sv"
`include "axi4_lite_scoreboard.sv"
`include "axi4_lite_env.sv"


endpackage 

//------------------------------------------------------------------------------------------------------------


